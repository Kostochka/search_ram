//////////////////////////////////////////////////////
// Module name:		parser_package
// Description: 	
// Originator:  	KOSTOCHKIN
// Rev:		Rev1.0 
// Date:	13_11_2019
// Project: 10G 
//////////////////////////////////////////////////////	

`timescale 1ns / 1ps   

package test_pkg; 

	const logic [0:32][7:0] data_arr_bytes_0 = 
	{
		8'h05, 8'h78, 8'h00, 8'h0E, 8'h01, 8'h01, 8'hBC, 8'h01, 8'h03, 8'h02, 8'h2B, 8'h01, 8'h03, 8'h09, 8'h01, 8'h03, 
		8'h03, 8'h78, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 
		8'h00
	}; 
	
	const logic [0:32][7:0] data_arr_bytes_1 = 
	{
		8'h05, 8'h78, 8'h00, 8'h15, 8'h01, 8'h01, 8'h4D, 8'h01, 8'h03, 8'h01, 8'hBC, 8'h01, 8'h01, 8'hBC, 8'h01, 8'h03, 
		8'h02, 8'h2B, 8'h01, 8'h03, 8'h09, 8'h01, 8'h03, 8'h03, 8'h78, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 
		8'h00
	};

	const logic [0:32][7:0] data_arr_bytes_2 = 
	{
		8'h00, 8'h00, 8'h00, 8'h1C, 8'h01, 8'h00, 8'hDE, 8'h01, 8'h03, 8'h01, 8'h4D, 8'h01, 8'h02, 8'h2B, 8'h01, 8'h03, 
		8'h02, 8'h9A, 8'h01, 8'h02, 8'h9A, 8'h01, 8'h03, 8'h03, 8'h09, 8'h01, 8'h03, 8'h78, 8'h01, 8'h03, 8'h03, 8'hE7, 
		8'hFF
	}; 	
	
	const logic [0:44][7:0] data_arr_bytes_3 = 
	{
		8'h00, 8'h00, 8'h00, 8'h07, 8'h01, 8'h02, 8'h9a, 8'h01, 8'h03, 8'h03, 8'h09, 8'hff, 8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00
	};
	
	const logic [0:44][7:0] data_arr_bytes_4 = 
	{
		8'h00, 8'h00, 8'h00, 8'h0e, 8'h01, 8'h00, 8'hde, 8'h01, 8'h03, 8'h01, 8'h4d, 8'h01, 8'h02, 8'h2b, 8'h01, 8'h03,
		8'h02, 8'h9a, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
		8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00	
	};
	
	const logic [0:44][7:0] data_arr_bytes_5 = 
	{
		8'h00, 8'h00, 8'h00, 8'h15, 8'h01, 8'h00, 8'hde, 8'h01, 8'h03, 8'h01, 8'h4d, 8'h01, 8'h02, 8'h2b, 8'h01, 8'h03, 
		8'h02, 8'h9a, 8'h01, 8'h03, 8'h78, 8'h01, 8'h03, 8'h03, 8'he7, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 
		8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00	
	};
	
	const logic [0:44][7:0] data_arr_bytes_6 = 
	{
		8'h05, 8'h78, 8'h00, 8'h15, 8'h01, 8'h01, 8'h4d, 8'h01, 8'h03, 8'h01, 8'hbc, 8'h01, 8'h01, 8'hbc, 8'h01, 8'h03, 
		8'h02, 8'h2b, 8'h01, 8'h03, 8'h09, 8'h01, 8'h03, 8'h03, 8'h78, 8'h01, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 
		8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00	
	};
	
	const logic [0:44][7:0] data_arr_bytes_7 = 
	{
		8'h00, 8'h00, 8'h00, 8'h1c, 8'h01, 8'h00, 8'hde, 8'h01, 8'h03, 8'h01, 8'h4d, 8'h01, 8'h02, 8'h2b, 8'h01, 8'h03, 
		8'h02, 8'h9a, 8'h01, 8'h02, 8'h9a, 8'h01, 8'h03, 8'h03, 8'h09, 8'h01, 8'h03, 8'h78, 8'h01, 8'h03, 8'h03, 8'he7,
		8'hff, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00	
	};


	const logic [0:67][55:0] data_arr_words = 
   {56'h000000_00007000,  //C
   
    56'h000001_00000000,  //D0
	56'h000003_10000011,  //D1
	56'h000006_10000111,  //D2
	56'h00000D_11111111,  //D3
	56'h00000E_00001111,  //D4
	56'h000300_10001111,  //D5
	56'h005000_00111110,  //D6
	56'h100000_00011110,  //D7
	56'hFFFFFF_11111110, 
	56'hFFFFFF_11110111,
	56'hFFFFFF_11111110, 
	56'hFFFFFF_11011111, 
	56'hFFFFFF_10111111, 
	56'hFFFFFF_11101111,
	56'hFFFFFF_11111101, 
	56'hFFFFFF_01111111,
	
	56'h000000_E0007000,  //C

    56'h000002_00000000,  //D0
	56'h000004_10100011,  //D1
	56'h000007_10100111,  //D2
	56'h00000A_11111111,  //D3
	56'h00000B_10001111,  //D4
	56'h00000C_10001111,  //D5
	56'h005001_10111110,  //D6
	56'h100100_10011110,  //D7
	56'hFFFFFF_11111110, 
	56'hFFFFFF_11110111,
	56'hFFFFFF_11111110, 
	56'hFFFFFF_11011111, 
	56'hFFFFFF_10111111, 
	56'hFFFFFF_11101111,
	56'hFFFFFF_11111101, 
	56'hFFFFFF_01111111,

	56'h000010_C0017000,  //C

    56'h000020_03000000,  //D0
	56'h000030_88888888,  //D1
	56'h000040_10150111,  //D2
	56'h000050_0A0A0A0A,  //D3
	56'h000060_10001B11,  //D4
	56'h000070_10C01111,  //D5
	56'h000080_AAAAAAAA,  //D6
	56'h000090_BBBBBBBB,  //D7
	56'h0000A0_CCCCCCCC, 
	56'h0000B0_DDDDDDDD,
	56'h0000C0_EEEEEEEE, 
	56'h0FFFFF_FFFFFFFF, 
	56'hFFFFFF_10111111, 
	56'hFFFFFF_11101111,
	56'hFFFFFF_11111101, 
	56'hFFFFFF_01111111,  	   
	
	56'h000010_A0027000,  //C
	
	56'h000011_B3000000,  //D0
	56'h000022_B8888888,  //D1
	56'h000033_B0150111,  //D2
	56'h000044_BA0A0A0A,  //D3
	56'h000055_B0001B11,  //D4
	56'h000066_B0C01111,  //D5
	56'h000077_CCCCCAAA,  //D6
	56'h000088_EEBBBBBB,  //D7
	56'h000099_88888888, 
	56'h0000AA_11111111,
	56'h0000BB_22345556, 
	56'h0000CC_98765432, 
	56'h0000DD_ABCCCDAE, 
	56'h0000EE_01010707,
	56'h0000FF_33333333, 
	56'h000FFF_09990009};
	
endpackage